module vaza (input I11,I12,I21,I22,I32,I33, output V,E,F);

	assign V = ((~I11)&(~I21)) | ((~I11)&(~I32)) | ((~I21)&(I33)) | ((~I21)&(I22)&(~I32)) | ((~I11)&(I22)&(I33)) | ((I22)&(~I32)&(I33)) | ((I12)&(I22)&(~I32));
	assign E = ((I11)&(I12)&(~I21)&(~I22)&(~I32)) | ((I11)&(I12)&(~I22)&(~I32)&(I33)) | ((I11)&(I12)&(~I21)&(I32)&(~I33)) | ((I11)&(I12)&(I21)&(I22)&(I32)&(I33));
	assign F = ((~I11)&(I12)&(I22)) | ((I12)&(~I21)&(I22)) | ((I12)&(I21)&(I33)) | ((I12)&(I21)&(I32)) | ((I11)&(I22)&(I33)) | ((I11)&(I22)&(I32)) | ((I11)&(~I12)&(I21)) | ((I11)&(I21)&(~I22));
	
endmodule 